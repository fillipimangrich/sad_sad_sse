library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
entity sad64pixels is
   PORT (
       v1,v2 : IN std_logic_vector(511 DOWNTO 0);
       q : OUT std_logic_vector(13 DOWNTO 0));
end sad64pixels;

architecture arch of sad64pixels is
begin
  q(7 downto 0) <= std_logic_vector(abs(signed(v1(7 downto 0)) - signed(v2(7 downto 0))));
  q(15 downto 8) <= std_logic_vector(abs(signed(v1(15 downto 8)) - signed(v2(15 downto 8))));
  q(23 downto 16) <= std_logic_vector(abs(signed(v1(23 downto 16)) - signed(v2(23 downto 16))));
  q(31 downto 24) <= std_logic_vector(abs(signed(v1(31 downto 24)) - signed(v2(31 downto 24))));
  q(39 downto 32) <= std_logic_vector(abs(signed(v1(39 downto 32)) - signed(v2(39 downto 32))));
  q(47 downto 40) <= std_logic_vector(abs(signed(v1(47 downto 40)) - signed(v2(47 downto 40))));
  q(55 downto 48) <= std_logic_vector(abs(signed(v1(55 downto 48)) - signed(v2(55 downto 48))));
  q(63 downto 56) <= std_logic_vector(abs(signed(v1(63 downto 56)) - signed(v2(63 downto 56))));
  q(71 downto 64) <= std_logic_vector(abs(signed(v1(71 downto 64)) - signed(v2(71 downto 64))));
  q(79 downto 72) <= std_logic_vector(abs(signed(v1(79 downto 72)) - signed(v2(79 downto 72))));
  q(87 downto 80) <= std_logic_vector(abs(signed(v1(87 downto 80)) - signed(v2(87 downto 80))));
  q(95 downto 88) <= std_logic_vector(abs(signed(v1(95 downto 88)) - signed(v2(95 downto 88))));
  q(103 downto 96) <= std_logic_vector(abs(signed(v1(103 downto 96)) - signed(v2(103 downto 96))));
  q(111 downto 104) <= std_logic_vector(abs(signed(v1(111 downto 104)) - signed(v2(111 downto 104))));
  q(119 downto 112) <= std_logic_vector(abs(signed(v1(119 downto 112)) - signed(v2(119 downto 112))));
  q(127 downto 120) <= std_logic_vector(abs(signed(v1(127 downto 120)) - signed(v2(127 downto 120))));
  q(135 downto 128) <= std_logic_vector(abs(signed(v1(135 downto 128)) - signed(v2(135 downto 128))));
  q(143 downto 136) <= std_logic_vector(abs(signed(v1(143 downto 136)) - signed(v2(143 downto 136))));
  q(151 downto 144) <= std_logic_vector(abs(signed(v1(151 downto 144)) - signed(v2(151 downto 144))));
  q(159 downto 152) <= std_logic_vector(abs(signed(v1(159 downto 152)) - signed(v2(159 downto 152))));
  q(167 downto 160) <= std_logic_vector(abs(signed(v1(167 downto 160)) - signed(v2(167 downto 160))));
  q(175 downto 168) <= std_logic_vector(abs(signed(v1(175 downto 168)) - signed(v2(175 downto 168))));
  q(183 downto 176) <= std_logic_vector(abs(signed(v1(183 downto 176)) - signed(v2(183 downto 176))));
  q(191 downto 184) <= std_logic_vector(abs(signed(v1(191 downto 184)) - signed(v2(191 downto 184))));
  q(199 downto 192) <= std_logic_vector(abs(signed(v1(199 downto 192)) - signed(v2(199 downto 192))));
  q(207 downto 200) <= std_logic_vector(abs(signed(v1(207 downto 200)) - signed(v2(207 downto 200))));
  q(215 downto 208) <= std_logic_vector(abs(signed(v1(215 downto 208)) - signed(v2(215 downto 208))));
  q(223 downto 216) <= std_logic_vector(abs(signed(v1(223 downto 216)) - signed(v2(223 downto 216))));
  q(231 downto 224) <= std_logic_vector(abs(signed(v1(231 downto 224)) - signed(v2(231 downto 224))));
  q(239 downto 232) <= std_logic_vector(abs(signed(v1(239 downto 232)) - signed(v2(239 downto 232))));
  q(247 downto 240) <= std_logic_vector(abs(signed(v1(247 downto 240)) - signed(v2(247 downto 240))));
  q(255 downto 248) <= std_logic_vector(abs(signed(v1(255 downto 248)) - signed(v2(255 downto 248))));
  q(263 downto 256) <= std_logic_vector(abs(signed(v1(263 downto 256)) - signed(v2(263 downto 256))));
  q(271 downto 264) <= std_logic_vector(abs(signed(v1(271 downto 264)) - signed(v2(271 downto 264))));
  q(279 downto 272) <= std_logic_vector(abs(signed(v1(279 downto 272)) - signed(v2(279 downto 272))));
  q(287 downto 280) <= std_logic_vector(abs(signed(v1(287 downto 280)) - signed(v2(287 downto 280))));
  q(295 downto 288) <= std_logic_vector(abs(signed(v1(295 downto 288)) - signed(v2(295 downto 288))));
  q(303 downto 296) <= std_logic_vector(abs(signed(v1(303 downto 296)) - signed(v2(303 downto 296))));
  q(311 downto 304) <= std_logic_vector(abs(signed(v1(311 downto 304)) - signed(v2(311 downto 304))));
  q(319 downto 312) <= std_logic_vector(abs(signed(v1(319 downto 312)) - signed(v2(319 downto 312))));
  q(327 downto 320) <= std_logic_vector(abs(signed(v1(327 downto 320)) - signed(v2(327 downto 320))));
  q(335 downto 328) <= std_logic_vector(abs(signed(v1(335 downto 328)) - signed(v2(335 downto 328))));
  q(343 downto 336) <= std_logic_vector(abs(signed(v1(343 downto 336)) - signed(v2(343 downto 336))));
  q(351 downto 344) <= std_logic_vector(abs(signed(v1(351 downto 344)) - signed(v2(351 downto 344))));
  q(359 downto 352) <= std_logic_vector(abs(signed(v1(359 downto 352)) - signed(v2(359 downto 352))));
  q(367 downto 360) <= std_logic_vector(abs(signed(v1(367 downto 360)) - signed(v2(367 downto 360))));
  q(375 downto 368) <= std_logic_vector(abs(signed(v1(375 downto 368)) - signed(v2(375 downto 368))));
  q(383 downto 376) <= std_logic_vector(abs(signed(v1(383 downto 376)) - signed(v2(383 downto 376))));
  q(391 downto 384) <= std_logic_vector(abs(signed(v1(391 downto 384)) - signed(v2(391 downto 384))));
  q(399 downto 392) <= std_logic_vector(abs(signed(v1(399 downto 392)) - signed(v2(399 downto 392))));
  q(407 downto 400) <= std_logic_vector(abs(signed(v1(407 downto 400)) - signed(v2(407 downto 400))));
  q(415 downto 408) <= std_logic_vector(abs(signed(v1(415 downto 408)) - signed(v2(415 downto 408))));
  q(423 downto 416) <= std_logic_vector(abs(signed(v1(423 downto 416)) - signed(v2(423 downto 416))));
  q(431 downto 424) <= std_logic_vector(abs(signed(v1(431 downto 424)) - signed(v2(431 downto 424))));
  q(439 downto 432) <= std_logic_vector(abs(signed(v1(439 downto 432)) - signed(v2(439 downto 432))));
  q(447 downto 440) <= std_logic_vector(abs(signed(v1(447 downto 440)) - signed(v2(447 downto 440))));
  q(455 downto 448) <= std_logic_vector(abs(signed(v1(455 downto 448)) - signed(v2(455 downto 448))));
  q(463 downto 456) <= std_logic_vector(abs(signed(v1(463 downto 456)) - signed(v2(463 downto 456))));
  q(471 downto 464) <= std_logic_vector(abs(signed(v1(471 downto 464)) - signed(v2(471 downto 464))));
  q(479 downto 472) <= std_logic_vector(abs(signed(v1(479 downto 472)) - signed(v2(479 downto 472))));
  q(487 downto 480) <= std_logic_vector(abs(signed(v1(487 downto 480)) - signed(v2(487 downto 480))));
  q(495 downto 488) <= std_logic_vector(abs(signed(v1(495 downto 488)) - signed(v2(495 downto 488))));
  q(503 downto 496) <= std_logic_vector(abs(signed(v1(503 downto 496)) - signed(v2(503 downto 496))));
  q(511 downto 504) <= std_logic_vector(abs(signed(v1(511 downto 504)) - signed(v2(511 downto 504))));
end arch;