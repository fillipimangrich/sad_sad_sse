library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity sum_tree_ssd128pixels is
   PORT (clk, enb, rst : IN STD_LOGIC;
       d : IN std_logic_vector(2047 DOWNTO 0);
       q : OUT std_logic_vector(22 DOWNTO 0));
end sum_tree_ssd128pixels;

architecture arch of sum_tree_ssd128pixels is
signal reg1, reg2, reg3, reg4, reg5, reg6, reg7, reg8, reg9, reg10, reg11, reg12, reg13, reg14, reg15, reg16, reg17, reg18, reg19, reg20, reg21, reg22, reg23, reg24, reg25, reg26, reg27, reg28, reg29, reg30, reg31, reg32, reg33, reg34, reg35, reg36, reg37, reg38, reg39, reg40, reg41, reg42, reg43, reg44, reg45, reg46, reg47, reg48, reg49, reg50, reg51, reg52, reg53, reg54, reg55, reg56, reg57, reg58, reg59, reg60, reg61, reg62, reg63, reg64 : std_logic_vector(16 downto 0);
signal reg65, reg66, reg67, reg68, reg69, reg70, reg71, reg72, reg73, reg74, reg75, reg76, reg77, reg78, reg79, reg80, reg81, reg82, reg83, reg84, reg85, reg86, reg87, reg88, reg89, reg90, reg91, reg92, reg93, reg94, reg95, reg96 : std_logic_vector(17 downto 0);
signal reg97, reg98, reg99, reg100, reg101, reg102, reg103, reg104, reg105, reg106, reg107, reg108, reg109, reg110, reg111, reg112 : std_logic_vector(18 downto 0);
signal reg113, reg114, reg115, reg116, reg117, reg118, reg119, reg120 : std_logic_vector(19 downto 0);
signal reg121, reg122, reg123, reg124 : std_logic_vector(20 downto 0);
signal reg125, reg126 : std_logic_vector(21 downto 0);
signal reg127 : std_logic_vector(22 downto 0);
BEGIN
   PROCESS(clk)
   BEGIN

       IF (rst = '1')THEN
           q <= (others => '0');
           reg1 <= (others => '0');
           reg2 <= (others => '0');
           reg3 <= (others => '0');
           reg4 <= (others => '0');
           reg5 <= (others => '0');
           reg6 <= (others => '0');
           reg7 <= (others => '0');
           reg8 <= (others => '0');
           reg9 <= (others => '0');
           reg10 <= (others => '0');
           reg11 <= (others => '0');
           reg12 <= (others => '0');
           reg13 <= (others => '0');
           reg14 <= (others => '0');
           reg15 <= (others => '0');
           reg16 <= (others => '0');
           reg17 <= (others => '0');
           reg18 <= (others => '0');
           reg19 <= (others => '0');
           reg20 <= (others => '0');
           reg21 <= (others => '0');
           reg22 <= (others => '0');
           reg23 <= (others => '0');
           reg24 <= (others => '0');
           reg25 <= (others => '0');
           reg26 <= (others => '0');
           reg27 <= (others => '0');
           reg28 <= (others => '0');
           reg29 <= (others => '0');
           reg30 <= (others => '0');
           reg31 <= (others => '0');
           reg32 <= (others => '0');
           reg33 <= (others => '0');
           reg34 <= (others => '0');
           reg35 <= (others => '0');
           reg36 <= (others => '0');
           reg37 <= (others => '0');
           reg38 <= (others => '0');
           reg39 <= (others => '0');
           reg40 <= (others => '0');
           reg41 <= (others => '0');
           reg42 <= (others => '0');
           reg43 <= (others => '0');
           reg44 <= (others => '0');
           reg45 <= (others => '0');
           reg46 <= (others => '0');
           reg47 <= (others => '0');
           reg48 <= (others => '0');
           reg49 <= (others => '0');
           reg50 <= (others => '0');
           reg51 <= (others => '0');
           reg52 <= (others => '0');
           reg53 <= (others => '0');
           reg54 <= (others => '0');
           reg55 <= (others => '0');
           reg56 <= (others => '0');
           reg57 <= (others => '0');
           reg58 <= (others => '0');
           reg59 <= (others => '0');
           reg60 <= (others => '0');
           reg61 <= (others => '0');
           reg62 <= (others => '0');
           reg63 <= (others => '0');
           reg64 <= (others => '0');
           reg65 <= (others => '0');
           reg66 <= (others => '0');
           reg67 <= (others => '0');
           reg68 <= (others => '0');
           reg69 <= (others => '0');
           reg70 <= (others => '0');
           reg71 <= (others => '0');
           reg72 <= (others => '0');
           reg73 <= (others => '0');
           reg74 <= (others => '0');
           reg75 <= (others => '0');
           reg76 <= (others => '0');
           reg77 <= (others => '0');
           reg78 <= (others => '0');
           reg79 <= (others => '0');
           reg80 <= (others => '0');
           reg81 <= (others => '0');
           reg82 <= (others => '0');
           reg83 <= (others => '0');
           reg84 <= (others => '0');
           reg85 <= (others => '0');
           reg86 <= (others => '0');
           reg87 <= (others => '0');
           reg88 <= (others => '0');
           reg89 <= (others => '0');
           reg90 <= (others => '0');
           reg91 <= (others => '0');
           reg92 <= (others => '0');
           reg93 <= (others => '0');
           reg94 <= (others => '0');
           reg95 <= (others => '0');
           reg96 <= (others => '0');
           reg97 <= (others => '0');
           reg98 <= (others => '0');
           reg99 <= (others => '0');
           reg100 <= (others => '0');
           reg101 <= (others => '0');
           reg102 <= (others => '0');
           reg103 <= (others => '0');
           reg104 <= (others => '0');
           reg105 <= (others => '0');
           reg106 <= (others => '0');
           reg107 <= (others => '0');
           reg108 <= (others => '0');
           reg109 <= (others => '0');
           reg110 <= (others => '0');
           reg111 <= (others => '0');
           reg112 <= (others => '0');
           reg113 <= (others => '0');
           reg114 <= (others => '0');
           reg115 <= (others => '0');
           reg116 <= (others => '0');
           reg117 <= (others => '0');
           reg118 <= (others => '0');
           reg119 <= (others => '0');
           reg120 <= (others => '0');
           reg121 <= (others => '0');
           reg122 <= (others => '0');
           reg123 <= (others => '0');
           reg124 <= (others => '0');
           reg125 <= (others => '0');
           reg126 <= (others => '0');
           reg127 <= (others => '0');
       ELSIF (clk'EVENT AND clk = '1' AND enb = '1') THEN
            reg1 <= ('0'&d(31 downto 16)) + ('0'&d(15 downto 0));
            reg2 <= ('0'&d(63 downto 48)) + ('0'&d(47 downto 32));
            reg3 <= ('0'&d(95 downto 80)) + ('0'&d(79 downto 64));
            reg4 <= ('0'&d(127 downto 112)) + ('0'&d(111 downto 96));
            reg5 <= ('0'&d(159 downto 144)) + ('0'&d(143 downto 128));
            reg6 <= ('0'&d(191 downto 176)) + ('0'&d(175 downto 160));
            reg7 <= ('0'&d(223 downto 208)) + ('0'&d(207 downto 192));
            reg8 <= ('0'&d(255 downto 240)) + ('0'&d(239 downto 224));
            reg9 <= ('0'&d(287 downto 272)) + ('0'&d(271 downto 256));
            reg10 <= ('0'&d(319 downto 304)) + ('0'&d(303 downto 288));
            reg11 <= ('0'&d(351 downto 336)) + ('0'&d(335 downto 320));
            reg12 <= ('0'&d(383 downto 368)) + ('0'&d(367 downto 352));
            reg13 <= ('0'&d(415 downto 400)) + ('0'&d(399 downto 384));
            reg14 <= ('0'&d(447 downto 432)) + ('0'&d(431 downto 416));
            reg15 <= ('0'&d(479 downto 464)) + ('0'&d(463 downto 448));
            reg16 <= ('0'&d(511 downto 496)) + ('0'&d(495 downto 480));
            reg17 <= ('0'&d(543 downto 528)) + ('0'&d(527 downto 512));
            reg18 <= ('0'&d(575 downto 560)) + ('0'&d(559 downto 544));
            reg19 <= ('0'&d(607 downto 592)) + ('0'&d(591 downto 576));
            reg20 <= ('0'&d(639 downto 624)) + ('0'&d(623 downto 608));
            reg21 <= ('0'&d(671 downto 656)) + ('0'&d(655 downto 640));
            reg22 <= ('0'&d(703 downto 688)) + ('0'&d(687 downto 672));
            reg23 <= ('0'&d(735 downto 720)) + ('0'&d(719 downto 704));
            reg24 <= ('0'&d(767 downto 752)) + ('0'&d(751 downto 736));
            reg25 <= ('0'&d(799 downto 784)) + ('0'&d(783 downto 768));
            reg26 <= ('0'&d(831 downto 816)) + ('0'&d(815 downto 800));
            reg27 <= ('0'&d(863 downto 848)) + ('0'&d(847 downto 832));
            reg28 <= ('0'&d(895 downto 880)) + ('0'&d(879 downto 864));
            reg29 <= ('0'&d(927 downto 912)) + ('0'&d(911 downto 896));
            reg30 <= ('0'&d(959 downto 944)) + ('0'&d(943 downto 928));
            reg31 <= ('0'&d(991 downto 976)) + ('0'&d(975 downto 960));
            reg32 <= ('0'&d(1023 downto 1008)) + ('0'&d(1007 downto 992));
            reg33 <= ('0'&d(1055 downto 1040)) + ('0'&d(1039 downto 1024));
            reg34 <= ('0'&d(1087 downto 1072)) + ('0'&d(1071 downto 1056));
            reg35 <= ('0'&d(1119 downto 1104)) + ('0'&d(1103 downto 1088));
            reg36 <= ('0'&d(1151 downto 1136)) + ('0'&d(1135 downto 1120));
            reg37 <= ('0'&d(1183 downto 1168)) + ('0'&d(1167 downto 1152));
            reg38 <= ('0'&d(1215 downto 1200)) + ('0'&d(1199 downto 1184));
            reg39 <= ('0'&d(1247 downto 1232)) + ('0'&d(1231 downto 1216));
            reg40 <= ('0'&d(1279 downto 1264)) + ('0'&d(1263 downto 1248));
            reg41 <= ('0'&d(1311 downto 1296)) + ('0'&d(1295 downto 1280));
            reg42 <= ('0'&d(1343 downto 1328)) + ('0'&d(1327 downto 1312));
            reg43 <= ('0'&d(1375 downto 1360)) + ('0'&d(1359 downto 1344));
            reg44 <= ('0'&d(1407 downto 1392)) + ('0'&d(1391 downto 1376));
            reg45 <= ('0'&d(1439 downto 1424)) + ('0'&d(1423 downto 1408));
            reg46 <= ('0'&d(1471 downto 1456)) + ('0'&d(1455 downto 1440));
            reg47 <= ('0'&d(1503 downto 1488)) + ('0'&d(1487 downto 1472));
            reg48 <= ('0'&d(1535 downto 1520)) + ('0'&d(1519 downto 1504));
            reg49 <= ('0'&d(1567 downto 1552)) + ('0'&d(1551 downto 1536));
            reg50 <= ('0'&d(1599 downto 1584)) + ('0'&d(1583 downto 1568));
            reg51 <= ('0'&d(1631 downto 1616)) + ('0'&d(1615 downto 1600));
            reg52 <= ('0'&d(1663 downto 1648)) + ('0'&d(1647 downto 1632));
            reg53 <= ('0'&d(1695 downto 1680)) + ('0'&d(1679 downto 1664));
            reg54 <= ('0'&d(1727 downto 1712)) + ('0'&d(1711 downto 1696));
            reg55 <= ('0'&d(1759 downto 1744)) + ('0'&d(1743 downto 1728));
            reg56 <= ('0'&d(1791 downto 1776)) + ('0'&d(1775 downto 1760));
            reg57 <= ('0'&d(1823 downto 1808)) + ('0'&d(1807 downto 1792));
            reg58 <= ('0'&d(1855 downto 1840)) + ('0'&d(1839 downto 1824));
            reg59 <= ('0'&d(1887 downto 1872)) + ('0'&d(1871 downto 1856));
            reg60 <= ('0'&d(1919 downto 1904)) + ('0'&d(1903 downto 1888));
            reg61 <= ('0'&d(1951 downto 1936)) + ('0'&d(1935 downto 1920));
            reg62 <= ('0'&d(1983 downto 1968)) + ('0'&d(1967 downto 1952));
            reg63 <= ('0'&d(2015 downto 2000)) + ('0'&d(1999 downto 1984));
            reg64 <= ('0'&d(2047 downto 2032)) + ('0'&d(2031 downto 2016));
            reg65 <= ('0'&reg1) + ('0'&reg2);
            reg66 <= ('0'&reg3) + ('0'&reg4);
            reg67 <= ('0'&reg5) + ('0'&reg6);
            reg68 <= ('0'&reg7) + ('0'&reg8);
            reg69 <= ('0'&reg9) + ('0'&reg10);
            reg70 <= ('0'&reg11) + ('0'&reg12);
            reg71 <= ('0'&reg13) + ('0'&reg14);
            reg72 <= ('0'&reg15) + ('0'&reg16);
            reg73 <= ('0'&reg17) + ('0'&reg18);
            reg74 <= ('0'&reg19) + ('0'&reg20);
            reg75 <= ('0'&reg21) + ('0'&reg22);
            reg76 <= ('0'&reg23) + ('0'&reg24);
            reg77 <= ('0'&reg25) + ('0'&reg26);
            reg78 <= ('0'&reg27) + ('0'&reg28);
            reg79 <= ('0'&reg29) + ('0'&reg30);
            reg80 <= ('0'&reg31) + ('0'&reg32);
            reg81 <= ('0'&reg33) + ('0'&reg34);
            reg82 <= ('0'&reg35) + ('0'&reg36);
            reg83 <= ('0'&reg37) + ('0'&reg38);
            reg84 <= ('0'&reg39) + ('0'&reg40);
            reg85 <= ('0'&reg41) + ('0'&reg42);
            reg86 <= ('0'&reg43) + ('0'&reg44);
            reg87 <= ('0'&reg45) + ('0'&reg46);
            reg88 <= ('0'&reg47) + ('0'&reg48);
            reg89 <= ('0'&reg49) + ('0'&reg50);
            reg90 <= ('0'&reg51) + ('0'&reg52);
            reg91 <= ('0'&reg53) + ('0'&reg54);
            reg92 <= ('0'&reg55) + ('0'&reg56);
            reg93 <= ('0'&reg57) + ('0'&reg58);
            reg94 <= ('0'&reg59) + ('0'&reg60);
            reg95 <= ('0'&reg61) + ('0'&reg62);
            reg96 <= ('0'&reg63) + ('0'&reg64);
            reg97 <= ('0'&reg65) + ('0'&reg66);
            reg98 <= ('0'&reg67) + ('0'&reg68);
            reg99 <= ('0'&reg69) + ('0'&reg70);
            reg100 <= ('0'&reg71) + ('0'&reg72);
            reg101 <= ('0'&reg73) + ('0'&reg74);
            reg102 <= ('0'&reg75) + ('0'&reg76);
            reg103 <= ('0'&reg77) + ('0'&reg78);
            reg104 <= ('0'&reg79) + ('0'&reg80);
            reg105 <= ('0'&reg81) + ('0'&reg82);
            reg106 <= ('0'&reg83) + ('0'&reg84);
            reg107 <= ('0'&reg85) + ('0'&reg86);
            reg108 <= ('0'&reg87) + ('0'&reg88);
            reg109 <= ('0'&reg89) + ('0'&reg90);
            reg110 <= ('0'&reg91) + ('0'&reg92);
            reg111 <= ('0'&reg93) + ('0'&reg94);
            reg112 <= ('0'&reg95) + ('0'&reg96);
            reg113 <= ('0'&reg97) + ('0'&reg98);
            reg114 <= ('0'&reg99) + ('0'&reg100);
            reg115 <= ('0'&reg101) + ('0'&reg102);
            reg116 <= ('0'&reg103) + ('0'&reg104);
            reg117 <= ('0'&reg105) + ('0'&reg106);
            reg118 <= ('0'&reg107) + ('0'&reg108);
            reg119 <= ('0'&reg109) + ('0'&reg110);
            reg120 <= ('0'&reg111) + ('0'&reg112);
            reg121 <= ('0'&reg113) + ('0'&reg114);
            reg122 <= ('0'&reg115) + ('0'&reg116);
            reg123 <= ('0'&reg117) + ('0'&reg118);
            reg124 <= ('0'&reg119) + ('0'&reg120);
            reg125 <= ('0'&reg121) + ('0'&reg122);
            reg126 <= ('0'&reg123) + ('0'&reg124);
            reg127 <= reg127 + ('0'&reg125) + ('0'&reg126);
        END IF;
          q <= reg127;
	END PROCESS;
END arch;