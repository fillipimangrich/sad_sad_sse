library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity sad16pixels is
   PORT (
       v1,v2 : IN std_logic_vector(127 DOWNTO 0);
       q : OUT std_logic_vector(127 DOWNTO 0));
end sad16pixels;

architecture arch of sad16pixels is
begin
  q(7 downto 0) <= std_logic_vector(abs(signed(v1(7 downto 0)) - signed(v2(7 downto 0))));
  q(15 downto 8) <= std_logic_vector(abs(signed(v1(15 downto 8)) - signed(v2(15 downto 8))));
  q(23 downto 16) <= std_logic_vector(abs(signed(v1(23 downto 16)) - signed(v2(23 downto 16))));
  q(31 downto 24) <= std_logic_vector(abs(signed(v1(31 downto 24)) - signed(v2(31 downto 24))));
  q(39 downto 32) <= std_logic_vector(abs(signed(v1(39 downto 32)) - signed(v2(39 downto 32))));
  q(47 downto 40) <= std_logic_vector(abs(signed(v1(47 downto 40)) - signed(v2(47 downto 40))));
  q(55 downto 48) <= std_logic_vector(abs(signed(v1(55 downto 48)) - signed(v2(55 downto 48))));
  q(63 downto 56) <= std_logic_vector(abs(signed(v1(63 downto 56)) - signed(v2(63 downto 56))));
  q(71 downto 64) <= std_logic_vector(abs(signed(v1(71 downto 64)) - signed(v2(71 downto 64))));
  q(79 downto 72) <= std_logic_vector(abs(signed(v1(79 downto 72)) - signed(v2(79 downto 72))));
  q(87 downto 80) <= std_logic_vector(abs(signed(v1(87 downto 80)) - signed(v2(87 downto 80))));
  q(95 downto 88) <= std_logic_vector(abs(signed(v1(95 downto 88)) - signed(v2(95 downto 88))));
  q(103 downto 96) <= std_logic_vector(abs(signed(v1(103 downto 96)) - signed(v2(103 downto 96))));
  q(111 downto 104) <= std_logic_vector(abs(signed(v1(111 downto 104)) - signed(v2(111 downto 104))));
  q(119 downto 112) <= std_logic_vector(abs(signed(v1(119 downto 112)) - signed(v2(119 downto 112))));
  q(127 downto 120) <= std_logic_vector(abs(signed(v1(127 downto 120)) - signed(v2(127 downto 120))));
end arch;