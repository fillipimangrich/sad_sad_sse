library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity sum_tree128pixels is
   PORT (clk, enb, rst : IN STD_LOGIC;
       d : IN std_logic_vector(1023 DOWNTO 0);
       q : OUT std_logic_vector(14 DOWNTO 0));
end sum_tree128pixels;

architecture arch of sum_tree128pixels is
signal reg1, reg2, reg3, reg4, reg5, reg6, reg7, reg8, reg9, reg10, reg11, reg12, reg13, reg14, reg15, reg16, reg17, reg18, reg19, reg20, reg21, reg22, reg23, reg24, reg25, reg26, reg27, reg28, reg29, reg30, reg31, reg32, reg33, reg34, reg35, reg36, reg37, reg38, reg39, reg40, reg41, reg42, reg43, reg44, reg45, reg46, reg47, reg48, reg49, reg50, reg51, reg52, reg53, reg54, reg55, reg56, reg57, reg58, reg59, reg60, reg61, reg62, reg63, reg64 : std_logic_vector(9 downto 0);
signal reg65, reg66, reg67, reg68, reg69, reg70, reg71, reg72, reg73, reg74, reg75, reg76, reg77, reg78, reg79, reg80, reg81, reg82, reg83, reg84, reg85, reg86, reg87, reg88, reg89, reg90, reg91, reg92, reg93, reg94, reg95, reg96 : std_logic_vector(10 downto 0);
signal reg97, reg98, reg99, reg100, reg101, reg102, reg103, reg104, reg105, reg106, reg107, reg108, reg109, reg110, reg111, reg112 : std_logic_vector(11 downto 0);
signal reg113, reg114, reg115, reg116, reg117, reg118, reg119, reg120 : std_logic_vector(12 downto 0);
signal reg121, reg122, reg123, reg124 : std_logic_vector(13 downto 0);
signal reg125, reg126 : std_logic_vector(14 downto 0);
signal reg127 : std_logic_vector(15 downto 0);
BEGIN
   PROCESS(clk)
   BEGIN

       IF (rst = 1)THEN
           q <= (others => '0');
           reg0 = (others => '0');
           reg1 = (others => '0');
           reg2 = (others => '0');
           reg3 = (others => '0');
           reg4 = (others => '0');
           reg5 = (others => '0');
           reg6 = (others => '0');
           reg7 = (others => '0');
           reg8 = (others => '0');
           reg9 = (others => '0');
           reg10 = (others => '0');
           reg11 = (others => '0');
           reg12 = (others => '0');
           reg13 = (others => '0');
           reg14 = (others => '0');
           reg15 = (others => '0');
           reg16 = (others => '0');
           reg17 = (others => '0');
           reg18 = (others => '0');
           reg19 = (others => '0');
           reg20 = (others => '0');
           reg21 = (others => '0');
           reg22 = (others => '0');
           reg23 = (others => '0');
           reg24 = (others => '0');
           reg25 = (others => '0');
           reg26 = (others => '0');
           reg27 = (others => '0');
           reg28 = (others => '0');
           reg29 = (others => '0');
           reg30 = (others => '0');
           reg31 = (others => '0');
           reg32 = (others => '0');
           reg33 = (others => '0');
           reg34 = (others => '0');
           reg35 = (others => '0');
           reg36 = (others => '0');
           reg37 = (others => '0');
           reg38 = (others => '0');
           reg39 = (others => '0');
           reg40 = (others => '0');
           reg41 = (others => '0');
           reg42 = (others => '0');
           reg43 = (others => '0');
           reg44 = (others => '0');
           reg45 = (others => '0');
           reg46 = (others => '0');
           reg47 = (others => '0');
           reg48 = (others => '0');
           reg49 = (others => '0');
           reg50 = (others => '0');
           reg51 = (others => '0');
           reg52 = (others => '0');
           reg53 = (others => '0');
           reg54 = (others => '0');
           reg55 = (others => '0');
           reg56 = (others => '0');
           reg57 = (others => '0');
           reg58 = (others => '0');
           reg59 = (others => '0');
           reg60 = (others => '0');
           reg61 = (others => '0');
           reg62 = (others => '0');
           reg63 = (others => '0');
           reg64 = (others => '0');
           reg65 = (others => '0');
           reg66 = (others => '0');
           reg67 = (others => '0');
           reg68 = (others => '0');
           reg69 = (others => '0');
           reg70 = (others => '0');
           reg71 = (others => '0');
           reg72 = (others => '0');
           reg73 = (others => '0');
           reg74 = (others => '0');
           reg75 = (others => '0');
           reg76 = (others => '0');
           reg77 = (others => '0');
           reg78 = (others => '0');
           reg79 = (others => '0');
           reg80 = (others => '0');
           reg81 = (others => '0');
           reg82 = (others => '0');
           reg83 = (others => '0');
           reg84 = (others => '0');
           reg85 = (others => '0');
           reg86 = (others => '0');
           reg87 = (others => '0');
           reg88 = (others => '0');
           reg89 = (others => '0');
           reg90 = (others => '0');
           reg91 = (others => '0');
           reg92 = (others => '0');
           reg93 = (others => '0');
           reg94 = (others => '0');
           reg95 = (others => '0');
           reg96 = (others => '0');
           reg97 = (others => '0');
           reg98 = (others => '0');
           reg99 = (others => '0');
           reg100 = (others => '0');
           reg101 = (others => '0');
           reg102 = (others => '0');
           reg103 = (others => '0');
           reg104 = (others => '0');
           reg105 = (others => '0');
           reg106 = (others => '0');
           reg107 = (others => '0');
           reg108 = (others => '0');
           reg109 = (others => '0');
           reg110 = (others => '0');
           reg111 = (others => '0');
           reg112 = (others => '0');
           reg113 = (others => '0');
           reg114 = (others => '0');
           reg115 = (others => '0');
           reg116 = (others => '0');
           reg117 = (others => '0');
           reg118 = (others => '0');
           reg119 = (others => '0');
           reg120 = (others => '0');
           reg121 = (others => '0');
           reg122 = (others => '0');
           reg123 = (others => '0');
           reg124 = (others => '0');
           reg125 = (others => '0');
           reg126 = (others => '0');
       ELSIF (clk'EVENT AND clk = '1' AND enb = '1') THEN
            reg1 <= ('0'&d(15 downto 8)) + ('0'&d(7 downto 0));
            reg2 <= ('0'&d(31 downto 24)) + ('0'&d(23 downto 16));
            reg3 <= ('0'&d(47 downto 40)) + ('0'&d(39 downto 32));
            reg4 <= ('0'&d(63 downto 56)) + ('0'&d(55 downto 48));
            reg5 <= ('0'&d(79 downto 72)) + ('0'&d(71 downto 64));
            reg6 <= ('0'&d(95 downto 88)) + ('0'&d(87 downto 80));
            reg7 <= ('0'&d(111 downto 104)) + ('0'&d(103 downto 96));
            reg8 <= ('0'&d(127 downto 120)) + ('0'&d(119 downto 112));
            reg9 <= ('0'&d(143 downto 136)) + ('0'&d(135 downto 128));
            reg10 <= ('0'&d(159 downto 152)) + ('0'&d(151 downto 144));
            reg11 <= ('0'&d(175 downto 168)) + ('0'&d(167 downto 160));
            reg12 <= ('0'&d(191 downto 184)) + ('0'&d(183 downto 176));
            reg13 <= ('0'&d(207 downto 200)) + ('0'&d(199 downto 192));
            reg14 <= ('0'&d(223 downto 216)) + ('0'&d(215 downto 208));
            reg15 <= ('0'&d(239 downto 232)) + ('0'&d(231 downto 224));
            reg16 <= ('0'&d(255 downto 248)) + ('0'&d(247 downto 240));
            reg17 <= ('0'&d(271 downto 264)) + ('0'&d(263 downto 256));
            reg18 <= ('0'&d(287 downto 280)) + ('0'&d(279 downto 272));
            reg19 <= ('0'&d(303 downto 296)) + ('0'&d(295 downto 288));
            reg20 <= ('0'&d(319 downto 312)) + ('0'&d(311 downto 304));
            reg21 <= ('0'&d(335 downto 328)) + ('0'&d(327 downto 320));
            reg22 <= ('0'&d(351 downto 344)) + ('0'&d(343 downto 336));
            reg23 <= ('0'&d(367 downto 360)) + ('0'&d(359 downto 352));
            reg24 <= ('0'&d(383 downto 376)) + ('0'&d(375 downto 368));
            reg25 <= ('0'&d(399 downto 392)) + ('0'&d(391 downto 384));
            reg26 <= ('0'&d(415 downto 408)) + ('0'&d(407 downto 400));
            reg27 <= ('0'&d(431 downto 424)) + ('0'&d(423 downto 416));
            reg28 <= ('0'&d(447 downto 440)) + ('0'&d(439 downto 432));
            reg29 <= ('0'&d(463 downto 456)) + ('0'&d(455 downto 448));
            reg30 <= ('0'&d(479 downto 472)) + ('0'&d(471 downto 464));
            reg31 <= ('0'&d(495 downto 488)) + ('0'&d(487 downto 480));
            reg32 <= ('0'&d(511 downto 504)) + ('0'&d(503 downto 496));
            reg33 <= ('0'&d(527 downto 520)) + ('0'&d(519 downto 512));
            reg34 <= ('0'&d(543 downto 536)) + ('0'&d(535 downto 528));
            reg35 <= ('0'&d(559 downto 552)) + ('0'&d(551 downto 544));
            reg36 <= ('0'&d(575 downto 568)) + ('0'&d(567 downto 560));
            reg37 <= ('0'&d(591 downto 584)) + ('0'&d(583 downto 576));
            reg38 <= ('0'&d(607 downto 600)) + ('0'&d(599 downto 592));
            reg39 <= ('0'&d(623 downto 616)) + ('0'&d(615 downto 608));
            reg40 <= ('0'&d(639 downto 632)) + ('0'&d(631 downto 624));
            reg41 <= ('0'&d(655 downto 648)) + ('0'&d(647 downto 640));
            reg42 <= ('0'&d(671 downto 664)) + ('0'&d(663 downto 656));
            reg43 <= ('0'&d(687 downto 680)) + ('0'&d(679 downto 672));
            reg44 <= ('0'&d(703 downto 696)) + ('0'&d(695 downto 688));
            reg45 <= ('0'&d(719 downto 712)) + ('0'&d(711 downto 704));
            reg46 <= ('0'&d(735 downto 728)) + ('0'&d(727 downto 720));
            reg47 <= ('0'&d(751 downto 744)) + ('0'&d(743 downto 736));
            reg48 <= ('0'&d(767 downto 760)) + ('0'&d(759 downto 752));
            reg49 <= ('0'&d(783 downto 776)) + ('0'&d(775 downto 768));
            reg50 <= ('0'&d(799 downto 792)) + ('0'&d(791 downto 784));
            reg51 <= ('0'&d(815 downto 808)) + ('0'&d(807 downto 800));
            reg52 <= ('0'&d(831 downto 824)) + ('0'&d(823 downto 816));
            reg53 <= ('0'&d(847 downto 840)) + ('0'&d(839 downto 832));
            reg54 <= ('0'&d(863 downto 856)) + ('0'&d(855 downto 848));
            reg55 <= ('0'&d(879 downto 872)) + ('0'&d(871 downto 864));
            reg56 <= ('0'&d(895 downto 888)) + ('0'&d(887 downto 880));
            reg57 <= ('0'&d(911 downto 904)) + ('0'&d(903 downto 896));
            reg58 <= ('0'&d(927 downto 920)) + ('0'&d(919 downto 912));
            reg59 <= ('0'&d(943 downto 936)) + ('0'&d(935 downto 928));
            reg60 <= ('0'&d(959 downto 952)) + ('0'&d(951 downto 944));
            reg61 <= ('0'&d(975 downto 968)) + ('0'&d(967 downto 960));
            reg62 <= ('0'&d(991 downto 984)) + ('0'&d(983 downto 976));
            reg63 <= ('0'&d(1007 downto 1000)) + ('0'&d(999 downto 992));
            reg64 <= ('0'&d(1023 downto 1016)) + ('0'&d(1015 downto 1008));
            reg65 <= ('0'&reg1) + ('0'&reg2);
            reg66 <= ('0'&reg3) + ('0'&reg4);
            reg67 <= ('0'&reg5) + ('0'&reg6);
            reg68 <= ('0'&reg7) + ('0'&reg8);
            reg69 <= ('0'&reg9) + ('0'&reg10);
            reg70 <= ('0'&reg11) + ('0'&reg12);
            reg71 <= ('0'&reg13) + ('0'&reg14);
            reg72 <= ('0'&reg15) + ('0'&reg16);
            reg73 <= ('0'&reg17) + ('0'&reg18);
            reg74 <= ('0'&reg19) + ('0'&reg20);
            reg75 <= ('0'&reg21) + ('0'&reg22);
            reg76 <= ('0'&reg23) + ('0'&reg24);
            reg77 <= ('0'&reg25) + ('0'&reg26);
            reg78 <= ('0'&reg27) + ('0'&reg28);
            reg79 <= ('0'&reg29) + ('0'&reg30);
            reg80 <= ('0'&reg31) + ('0'&reg32);
            reg81 <= ('0'&reg33) + ('0'&reg34);
            reg82 <= ('0'&reg35) + ('0'&reg36);
            reg83 <= ('0'&reg37) + ('0'&reg38);
            reg84 <= ('0'&reg39) + ('0'&reg40);
            reg85 <= ('0'&reg41) + ('0'&reg42);
            reg86 <= ('0'&reg43) + ('0'&reg44);
            reg87 <= ('0'&reg45) + ('0'&reg46);
            reg88 <= ('0'&reg47) + ('0'&reg48);
            reg89 <= ('0'&reg49) + ('0'&reg50);
            reg90 <= ('0'&reg51) + ('0'&reg52);
            reg91 <= ('0'&reg53) + ('0'&reg54);
            reg92 <= ('0'&reg55) + ('0'&reg56);
            reg93 <= ('0'&reg57) + ('0'&reg58);
            reg94 <= ('0'&reg59) + ('0'&reg60);
            reg95 <= ('0'&reg61) + ('0'&reg62);
            reg96 <= ('0'&reg63) + ('0'&reg64);
            reg97 <= ('0'&reg65) + ('0'&reg66);
            reg98 <= ('0'&reg67) + ('0'&reg68);
            reg99 <= ('0'&reg69) + ('0'&reg70);
            reg100 <= ('0'&reg71) + ('0'&reg72);
            reg101 <= ('0'&reg73) + ('0'&reg74);
            reg102 <= ('0'&reg75) + ('0'&reg76);
            reg103 <= ('0'&reg77) + ('0'&reg78);
            reg104 <= ('0'&reg79) + ('0'&reg80);
            reg105 <= ('0'&reg81) + ('0'&reg82);
            reg106 <= ('0'&reg83) + ('0'&reg84);
            reg107 <= ('0'&reg85) + ('0'&reg86);
            reg108 <= ('0'&reg87) + ('0'&reg88);
            reg109 <= ('0'&reg89) + ('0'&reg90);
            reg110 <= ('0'&reg91) + ('0'&reg92);
            reg111 <= ('0'&reg93) + ('0'&reg94);
            reg112 <= ('0'&reg95) + ('0'&reg96);
            reg113 <= ('0'&reg97) + ('0'&reg98);
            reg114 <= ('0'&reg99) + ('0'&reg100);
            reg115 <= ('0'&reg101) + ('0'&reg102);
            reg116 <= ('0'&reg103) + ('0'&reg104);
            reg117 <= ('0'&reg105) + ('0'&reg106);
            reg118 <= ('0'&reg107) + ('0'&reg108);
            reg119 <= ('0'&reg109) + ('0'&reg110);
            reg120 <= ('0'&reg111) + ('0'&reg112);
            reg121 <= ('0'&reg113) + ('0'&reg114);
            reg122 <= ('0'&reg115) + ('0'&reg116);
            reg123 <= ('0'&reg117) + ('0'&reg118);
            reg124 <= ('0'&reg119) + ('0'&reg120);
            reg125 <= ('0'&reg121) + ('0'&reg122);
            reg126 <= ('0'&reg123) + ('0'&reg124);
            reg127 <= reg127 + ('0'&reg125) + ('0'&reg126);
        END IF;
          q <= reg127;
	END PROCESS;
END arch;