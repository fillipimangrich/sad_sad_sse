library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity sum_tree is
   PORT (clk, enb, rst : IN STD_LOGIC;
       d : IN std_logic_vector(1023 DOWNTO 0);
       q : OUT std_logic_vector(21 DOWNTO 0));
end sum_tree;

architecture arch of sum_tree is
signal ZEROS : std_logic_vector(N - 1 DOWNTO 0) := (OTHERS => '0');
signal reg1, reg2, reg3, reg4, reg5, reg6, reg7, reg8, reg9, reg10, reg11, reg12, reg13, reg14, reg15, reg16, reg17, reg18, reg19, reg20, reg21, reg22, reg23, reg24, reg25, reg26, reg27, reg28, reg29, reg30, reg31, reg32, reg33, reg34, reg35, reg36, reg37, reg38, reg39, reg40, reg41, reg42, reg43, reg44, reg45, reg46, reg47, reg48, reg49, reg50, reg51, reg52, reg53, reg54, reg55, reg56, reg57, reg58, reg59, reg60, reg61, reg62, reg63, reg64 : std_logic_vector(129 downto 0);
signal reg65, reg66, reg67, reg68, reg69, reg70, reg71, reg72, reg73, reg74, reg75, reg76, reg77, reg78, reg79, reg80, reg81, reg82, reg83, reg84, reg85, reg86, reg87, reg88, reg89, reg90, reg91, reg92, reg93, reg94, reg95, reg96 : std_logic_vector(130 downto 0);
signal reg97, reg98, reg99, reg100, reg101, reg102, reg103, reg104, reg105, reg106, reg107, reg108, reg109, reg110, reg111, reg112, reg113, reg114, reg115, reg116, reg117 : std_logic_vector(131 downto 0);
signal reg118, reg119, reg120, reg121, reg122, reg123, reg124, reg125, reg126, reg127, reg128, reg129, reg130, reg131, reg132, reg133 : std_logic_vector(132 downto 0);
signal reg134, reg135, reg136, reg137, reg138, reg139, reg140, reg141, reg142, reg143, reg144, reg145 : std_logic_vector(133 downto 0);
signal reg146, reg147, reg148, reg149, reg150, reg151, reg152, reg153, reg154, reg155 : std_logic_vector(134 downto 0);
signal reg156, reg157, reg158, reg159, reg160, reg161, reg162, reg163, reg164 : std_logic_vector(135 downto 0);
BEGIN
   PROCESS(clk)
   BEGIN

       IF (rst = 1)THEN
           q <= (others => '0');
       ELSIF (clk'EVENT AND clk = '1' AND enb = '1') THEN
            reg1 <= '0'&d(15 downto 8) + '0'&d(7 downto 0);
            reg2 <= '0'&d(271 downto 264) + '0'&d(263 downto 256);
            reg3 <= '0'&d(527 downto 520) + '0'&d(519 downto 512);
            reg4 <= '0'&d(783 downto 776) + '0'&d(775 downto 768);
            reg5 <= '0'&d(1039 downto 1032) + '0'&d(1031 downto 1024);
            reg6 <= '0'&d(1295 downto 1288) + '0'&d(1287 downto 1280);
            reg7 <= '0'&d(1551 downto 1544) + '0'&d(1543 downto 1536);
            reg8 <= '0'&d(1807 downto 1800) + '0'&d(1799 downto 1792);
            reg9 <= '0'&d(2063 downto 2056) + '0'&d(2055 downto 2048);
            reg10 <= '0'&d(2319 downto 2312) + '0'&d(2311 downto 2304);
            reg11 <= '0'&d(2575 downto 2568) + '0'&d(2567 downto 2560);
            reg12 <= '0'&d(2831 downto 2824) + '0'&d(2823 downto 2816);
            reg13 <= '0'&d(3087 downto 3080) + '0'&d(3079 downto 3072);
            reg14 <= '0'&d(3343 downto 3336) + '0'&d(3335 downto 3328);
            reg15 <= '0'&d(3599 downto 3592) + '0'&d(3591 downto 3584);
            reg16 <= '0'&d(3855 downto 3848) + '0'&d(3847 downto 3840);
            reg17 <= '0'&d(4111 downto 4104) + '0'&d(4103 downto 4096);
            reg18 <= '0'&d(4367 downto 4360) + '0'&d(4359 downto 4352);
            reg19 <= '0'&d(4623 downto 4616) + '0'&d(4615 downto 4608);
            reg20 <= '0'&d(4879 downto 4872) + '0'&d(4871 downto 4864);
            reg21 <= '0'&d(5135 downto 5128) + '0'&d(5127 downto 5120);
            reg22 <= '0'&d(5391 downto 5384) + '0'&d(5383 downto 5376);
            reg23 <= '0'&d(5647 downto 5640) + '0'&d(5639 downto 5632);
            reg24 <= '0'&d(5903 downto 5896) + '0'&d(5895 downto 5888);
            reg25 <= '0'&d(6159 downto 6152) + '0'&d(6151 downto 6144);
            reg26 <= '0'&d(6415 downto 6408) + '0'&d(6407 downto 6400);
            reg27 <= '0'&d(6671 downto 6664) + '0'&d(6663 downto 6656);
            reg28 <= '0'&d(6927 downto 6920) + '0'&d(6919 downto 6912);
            reg29 <= '0'&d(7183 downto 7176) + '0'&d(7175 downto 7168);
            reg30 <= '0'&d(7439 downto 7432) + '0'&d(7431 downto 7424);
            reg31 <= '0'&d(7695 downto 7688) + '0'&d(7687 downto 7680);
            reg32 <= '0'&d(7951 downto 7944) + '0'&d(7943 downto 7936);
            reg33 <= '0'&d(8207 downto 8200) + '0'&d(8199 downto 8192);
            reg34 <= '0'&d(8463 downto 8456) + '0'&d(8455 downto 8448);
            reg35 <= '0'&d(8719 downto 8712) + '0'&d(8711 downto 8704);
            reg36 <= '0'&d(8975 downto 8968) + '0'&d(8967 downto 8960);
            reg37 <= '0'&d(9231 downto 9224) + '0'&d(9223 downto 9216);
            reg38 <= '0'&d(9487 downto 9480) + '0'&d(9479 downto 9472);
            reg39 <= '0'&d(9743 downto 9736) + '0'&d(9735 downto 9728);
            reg40 <= '0'&d(9999 downto 9992) + '0'&d(9991 downto 9984);
            reg41 <= '0'&d(10255 downto 10248) + '0'&d(10247 downto 10240);
            reg42 <= '0'&d(10511 downto 10504) + '0'&d(10503 downto 10496);
            reg43 <= '0'&d(10767 downto 10760) + '0'&d(10759 downto 10752);
            reg44 <= '0'&d(11023 downto 11016) + '0'&d(11015 downto 11008);
            reg45 <= '0'&d(11279 downto 11272) + '0'&d(11271 downto 11264);
            reg46 <= '0'&d(11535 downto 11528) + '0'&d(11527 downto 11520);
            reg47 <= '0'&d(11791 downto 11784) + '0'&d(11783 downto 11776);
            reg48 <= '0'&d(12047 downto 12040) + '0'&d(12039 downto 12032);
            reg49 <= '0'&d(12303 downto 12296) + '0'&d(12295 downto 12288);
            reg50 <= '0'&d(12559 downto 12552) + '0'&d(12551 downto 12544);
            reg51 <= '0'&d(12815 downto 12808) + '0'&d(12807 downto 12800);
            reg52 <= '0'&d(13071 downto 13064) + '0'&d(13063 downto 13056);
            reg53 <= '0'&d(13327 downto 13320) + '0'&d(13319 downto 13312);
            reg54 <= '0'&d(13583 downto 13576) + '0'&d(13575 downto 13568);
            reg55 <= '0'&d(13839 downto 13832) + '0'&d(13831 downto 13824);
            reg56 <= '0'&d(14095 downto 14088) + '0'&d(14087 downto 14080);
            reg57 <= '0'&d(14351 downto 14344) + '0'&d(14343 downto 14336);
            reg58 <= '0'&d(14607 downto 14600) + '0'&d(14599 downto 14592);
            reg59 <= '0'&d(14863 downto 14856) + '0'&d(14855 downto 14848);
            reg60 <= '0'&d(15119 downto 15112) + '0'&d(15111 downto 15104);
            reg61 <= '0'&d(15375 downto 15368) + '0'&d(15367 downto 15360);
            reg62 <= '0'&d(15631 downto 15624) + '0'&d(15623 downto 15616);
            reg63 <= '0'&d(15887 downto 15880) + '0'&d(15879 downto 15872);
            reg64 <= '0'&d(16143 downto 16136) + '0'&d(16135 downto 16128);
            reg65 <= reg1 + reg2;
            reg66 <= reg3 + reg4;
            reg67 <= reg5 + reg6;
            reg68 <= reg7 + reg8;
            reg69 <= reg9 + reg10;
            reg70 <= reg11 + reg12;
            reg71 <= reg13 + reg14;
            reg72 <= reg15 + reg16;
            reg73 <= reg17 + reg18;
            reg74 <= reg19 + reg20;
            reg75 <= reg21 + reg22;
            reg76 <= reg23 + reg24;
            reg77 <= reg25 + reg26;
            reg78 <= reg27 + reg28;
            reg79 <= reg29 + reg30;
            reg80 <= reg31 + reg32;
            reg81 <= reg33 + reg34;
            reg82 <= reg35 + reg36;
            reg83 <= reg37 + reg38;
            reg84 <= reg39 + reg40;
            reg85 <= reg41 + reg42;
            reg86 <= reg43 + reg44;
            reg87 <= reg45 + reg46;
            reg88 <= reg47 + reg48;
            reg89 <= reg49 + reg50;
            reg90 <= reg51 + reg52;
            reg91 <= reg53 + reg54;
            reg92 <= reg55 + reg56;
            reg93 <= reg57 + reg58;
            reg94 <= reg59 + reg60;
            reg95 <= reg61 + reg62;
            reg96 <= reg63 + reg64;
            reg97 <= reg65 + reg66;
            reg98 <= reg67 + reg68;
            reg99 <= reg69 + reg70;
            reg100 <= reg71 + reg72;
            reg101 <= reg73 + reg74;
            reg102 <= reg75 + reg76;
            reg103 <= reg77 + reg78;
            reg104 <= reg79 + reg80;
            reg105 <= reg81 + reg82;
            reg106 <= reg83 + reg84;
            reg107 <= reg85 + reg86;
            reg108 <= reg87 + reg88;
            reg109 <= reg89 + reg90;
            reg110 <= reg91 + reg92;
            reg111 <= reg93 + reg94;
            reg112 <= reg95 + reg96;
            reg113 <= reg97 + reg98;
            reg114 <= reg99 + reg100;
            reg115 <= reg101 + reg102;
            reg116 <= reg103 + reg104;
            reg117 <= reg105 + reg106;
            reg118 <= reg107 + reg108;
            reg119 <= reg109 + reg110;
            reg120 <= reg111 + reg112;
            reg121 <= reg113 + reg114;
            reg122 <= reg115 + reg116;
            reg123 <= reg117 + reg118;
            reg124 <= reg119 + reg120;
            reg125 <= reg121 + reg122;
            reg126 <= reg123 + reg124;
            reg127 <= reg127 + reg125 + reg126;
        END IF;
	END PROCESS;
q <= reg127;
END arch;