library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
entity sad128pixels is
   PORT (
       v1,v2 : IN std_logic_vector(1023 DOWNTO 0);
       q : OUT std_logic_vector(1023 DOWNTO 0));
end sad128pixels;

architecture arch of sad128pixels is
begin
  q(7 downto 0) <= std_logic_vector(abs(signed(v1(7 downto 0)) - signed(v2(7 downto 0))));
  q(15 downto 8) <= std_logic_vector(abs(signed(v1(15 downto 8)) - signed(v2(15 downto 8))));
  q(23 downto 16) <= std_logic_vector(abs(signed(v1(23 downto 16)) - signed(v2(23 downto 16))));
  q(31 downto 24) <= std_logic_vector(abs(signed(v1(31 downto 24)) - signed(v2(31 downto 24))));
  q(39 downto 32) <= std_logic_vector(abs(signed(v1(39 downto 32)) - signed(v2(39 downto 32))));
  q(47 downto 40) <= std_logic_vector(abs(signed(v1(47 downto 40)) - signed(v2(47 downto 40))));
  q(55 downto 48) <= std_logic_vector(abs(signed(v1(55 downto 48)) - signed(v2(55 downto 48))));
  q(63 downto 56) <= std_logic_vector(abs(signed(v1(63 downto 56)) - signed(v2(63 downto 56))));
  q(71 downto 64) <= std_logic_vector(abs(signed(v1(71 downto 64)) - signed(v2(71 downto 64))));
  q(79 downto 72) <= std_logic_vector(abs(signed(v1(79 downto 72)) - signed(v2(79 downto 72))));
  q(87 downto 80) <= std_logic_vector(abs(signed(v1(87 downto 80)) - signed(v2(87 downto 80))));
  q(95 downto 88) <= std_logic_vector(abs(signed(v1(95 downto 88)) - signed(v2(95 downto 88))));
  q(103 downto 96) <= std_logic_vector(abs(signed(v1(103 downto 96)) - signed(v2(103 downto 96))));
  q(111 downto 104) <= std_logic_vector(abs(signed(v1(111 downto 104)) - signed(v2(111 downto 104))));
  q(119 downto 112) <= std_logic_vector(abs(signed(v1(119 downto 112)) - signed(v2(119 downto 112))));
  q(127 downto 120) <= std_logic_vector(abs(signed(v1(127 downto 120)) - signed(v2(127 downto 120))));
  q(135 downto 128) <= std_logic_vector(abs(signed(v1(135 downto 128)) - signed(v2(135 downto 128))));
  q(143 downto 136) <= std_logic_vector(abs(signed(v1(143 downto 136)) - signed(v2(143 downto 136))));
  q(151 downto 144) <= std_logic_vector(abs(signed(v1(151 downto 144)) - signed(v2(151 downto 144))));
  q(159 downto 152) <= std_logic_vector(abs(signed(v1(159 downto 152)) - signed(v2(159 downto 152))));
  q(167 downto 160) <= std_logic_vector(abs(signed(v1(167 downto 160)) - signed(v2(167 downto 160))));
  q(175 downto 168) <= std_logic_vector(abs(signed(v1(175 downto 168)) - signed(v2(175 downto 168))));
  q(183 downto 176) <= std_logic_vector(abs(signed(v1(183 downto 176)) - signed(v2(183 downto 176))));
  q(191 downto 184) <= std_logic_vector(abs(signed(v1(191 downto 184)) - signed(v2(191 downto 184))));
  q(199 downto 192) <= std_logic_vector(abs(signed(v1(199 downto 192)) - signed(v2(199 downto 192))));
  q(207 downto 200) <= std_logic_vector(abs(signed(v1(207 downto 200)) - signed(v2(207 downto 200))));
  q(215 downto 208) <= std_logic_vector(abs(signed(v1(215 downto 208)) - signed(v2(215 downto 208))));
  q(223 downto 216) <= std_logic_vector(abs(signed(v1(223 downto 216)) - signed(v2(223 downto 216))));
  q(231 downto 224) <= std_logic_vector(abs(signed(v1(231 downto 224)) - signed(v2(231 downto 224))));
  q(239 downto 232) <= std_logic_vector(abs(signed(v1(239 downto 232)) - signed(v2(239 downto 232))));
  q(247 downto 240) <= std_logic_vector(abs(signed(v1(247 downto 240)) - signed(v2(247 downto 240))));
  q(255 downto 248) <= std_logic_vector(abs(signed(v1(255 downto 248)) - signed(v2(255 downto 248))));
  q(263 downto 256) <= std_logic_vector(abs(signed(v1(263 downto 256)) - signed(v2(263 downto 256))));
  q(271 downto 264) <= std_logic_vector(abs(signed(v1(271 downto 264)) - signed(v2(271 downto 264))));
  q(279 downto 272) <= std_logic_vector(abs(signed(v1(279 downto 272)) - signed(v2(279 downto 272))));
  q(287 downto 280) <= std_logic_vector(abs(signed(v1(287 downto 280)) - signed(v2(287 downto 280))));
  q(295 downto 288) <= std_logic_vector(abs(signed(v1(295 downto 288)) - signed(v2(295 downto 288))));
  q(303 downto 296) <= std_logic_vector(abs(signed(v1(303 downto 296)) - signed(v2(303 downto 296))));
  q(311 downto 304) <= std_logic_vector(abs(signed(v1(311 downto 304)) - signed(v2(311 downto 304))));
  q(319 downto 312) <= std_logic_vector(abs(signed(v1(319 downto 312)) - signed(v2(319 downto 312))));
  q(327 downto 320) <= std_logic_vector(abs(signed(v1(327 downto 320)) - signed(v2(327 downto 320))));
  q(335 downto 328) <= std_logic_vector(abs(signed(v1(335 downto 328)) - signed(v2(335 downto 328))));
  q(343 downto 336) <= std_logic_vector(abs(signed(v1(343 downto 336)) - signed(v2(343 downto 336))));
  q(351 downto 344) <= std_logic_vector(abs(signed(v1(351 downto 344)) - signed(v2(351 downto 344))));
  q(359 downto 352) <= std_logic_vector(abs(signed(v1(359 downto 352)) - signed(v2(359 downto 352))));
  q(367 downto 360) <= std_logic_vector(abs(signed(v1(367 downto 360)) - signed(v2(367 downto 360))));
  q(375 downto 368) <= std_logic_vector(abs(signed(v1(375 downto 368)) - signed(v2(375 downto 368))));
  q(383 downto 376) <= std_logic_vector(abs(signed(v1(383 downto 376)) - signed(v2(383 downto 376))));
  q(391 downto 384) <= std_logic_vector(abs(signed(v1(391 downto 384)) - signed(v2(391 downto 384))));
  q(399 downto 392) <= std_logic_vector(abs(signed(v1(399 downto 392)) - signed(v2(399 downto 392))));
  q(407 downto 400) <= std_logic_vector(abs(signed(v1(407 downto 400)) - signed(v2(407 downto 400))));
  q(415 downto 408) <= std_logic_vector(abs(signed(v1(415 downto 408)) - signed(v2(415 downto 408))));
  q(423 downto 416) <= std_logic_vector(abs(signed(v1(423 downto 416)) - signed(v2(423 downto 416))));
  q(431 downto 424) <= std_logic_vector(abs(signed(v1(431 downto 424)) - signed(v2(431 downto 424))));
  q(439 downto 432) <= std_logic_vector(abs(signed(v1(439 downto 432)) - signed(v2(439 downto 432))));
  q(447 downto 440) <= std_logic_vector(abs(signed(v1(447 downto 440)) - signed(v2(447 downto 440))));
  q(455 downto 448) <= std_logic_vector(abs(signed(v1(455 downto 448)) - signed(v2(455 downto 448))));
  q(463 downto 456) <= std_logic_vector(abs(signed(v1(463 downto 456)) - signed(v2(463 downto 456))));
  q(471 downto 464) <= std_logic_vector(abs(signed(v1(471 downto 464)) - signed(v2(471 downto 464))));
  q(479 downto 472) <= std_logic_vector(abs(signed(v1(479 downto 472)) - signed(v2(479 downto 472))));
  q(487 downto 480) <= std_logic_vector(abs(signed(v1(487 downto 480)) - signed(v2(487 downto 480))));
  q(495 downto 488) <= std_logic_vector(abs(signed(v1(495 downto 488)) - signed(v2(495 downto 488))));
  q(503 downto 496) <= std_logic_vector(abs(signed(v1(503 downto 496)) - signed(v2(503 downto 496))));
  q(511 downto 504) <= std_logic_vector(abs(signed(v1(511 downto 504)) - signed(v2(511 downto 504))));
  q(519 downto 512) <= std_logic_vector(abs(signed(v1(519 downto 512)) - signed(v2(519 downto 512))));
  q(527 downto 520) <= std_logic_vector(abs(signed(v1(527 downto 520)) - signed(v2(527 downto 520))));
  q(535 downto 528) <= std_logic_vector(abs(signed(v1(535 downto 528)) - signed(v2(535 downto 528))));
  q(543 downto 536) <= std_logic_vector(abs(signed(v1(543 downto 536)) - signed(v2(543 downto 536))));
  q(551 downto 544) <= std_logic_vector(abs(signed(v1(551 downto 544)) - signed(v2(551 downto 544))));
  q(559 downto 552) <= std_logic_vector(abs(signed(v1(559 downto 552)) - signed(v2(559 downto 552))));
  q(567 downto 560) <= std_logic_vector(abs(signed(v1(567 downto 560)) - signed(v2(567 downto 560))));
  q(575 downto 568) <= std_logic_vector(abs(signed(v1(575 downto 568)) - signed(v2(575 downto 568))));
  q(583 downto 576) <= std_logic_vector(abs(signed(v1(583 downto 576)) - signed(v2(583 downto 576))));
  q(591 downto 584) <= std_logic_vector(abs(signed(v1(591 downto 584)) - signed(v2(591 downto 584))));
  q(599 downto 592) <= std_logic_vector(abs(signed(v1(599 downto 592)) - signed(v2(599 downto 592))));
  q(607 downto 600) <= std_logic_vector(abs(signed(v1(607 downto 600)) - signed(v2(607 downto 600))));
  q(615 downto 608) <= std_logic_vector(abs(signed(v1(615 downto 608)) - signed(v2(615 downto 608))));
  q(623 downto 616) <= std_logic_vector(abs(signed(v1(623 downto 616)) - signed(v2(623 downto 616))));
  q(631 downto 624) <= std_logic_vector(abs(signed(v1(631 downto 624)) - signed(v2(631 downto 624))));
  q(639 downto 632) <= std_logic_vector(abs(signed(v1(639 downto 632)) - signed(v2(639 downto 632))));
  q(647 downto 640) <= std_logic_vector(abs(signed(v1(647 downto 640)) - signed(v2(647 downto 640))));
  q(655 downto 648) <= std_logic_vector(abs(signed(v1(655 downto 648)) - signed(v2(655 downto 648))));
  q(663 downto 656) <= std_logic_vector(abs(signed(v1(663 downto 656)) - signed(v2(663 downto 656))));
  q(671 downto 664) <= std_logic_vector(abs(signed(v1(671 downto 664)) - signed(v2(671 downto 664))));
  q(679 downto 672) <= std_logic_vector(abs(signed(v1(679 downto 672)) - signed(v2(679 downto 672))));
  q(687 downto 680) <= std_logic_vector(abs(signed(v1(687 downto 680)) - signed(v2(687 downto 680))));
  q(695 downto 688) <= std_logic_vector(abs(signed(v1(695 downto 688)) - signed(v2(695 downto 688))));
  q(703 downto 696) <= std_logic_vector(abs(signed(v1(703 downto 696)) - signed(v2(703 downto 696))));
  q(711 downto 704) <= std_logic_vector(abs(signed(v1(711 downto 704)) - signed(v2(711 downto 704))));
  q(719 downto 712) <= std_logic_vector(abs(signed(v1(719 downto 712)) - signed(v2(719 downto 712))));
  q(727 downto 720) <= std_logic_vector(abs(signed(v1(727 downto 720)) - signed(v2(727 downto 720))));
  q(735 downto 728) <= std_logic_vector(abs(signed(v1(735 downto 728)) - signed(v2(735 downto 728))));
  q(743 downto 736) <= std_logic_vector(abs(signed(v1(743 downto 736)) - signed(v2(743 downto 736))));
  q(751 downto 744) <= std_logic_vector(abs(signed(v1(751 downto 744)) - signed(v2(751 downto 744))));
  q(759 downto 752) <= std_logic_vector(abs(signed(v1(759 downto 752)) - signed(v2(759 downto 752))));
  q(767 downto 760) <= std_logic_vector(abs(signed(v1(767 downto 760)) - signed(v2(767 downto 760))));
  q(775 downto 768) <= std_logic_vector(abs(signed(v1(775 downto 768)) - signed(v2(775 downto 768))));
  q(783 downto 776) <= std_logic_vector(abs(signed(v1(783 downto 776)) - signed(v2(783 downto 776))));
  q(791 downto 784) <= std_logic_vector(abs(signed(v1(791 downto 784)) - signed(v2(791 downto 784))));
  q(799 downto 792) <= std_logic_vector(abs(signed(v1(799 downto 792)) - signed(v2(799 downto 792))));
  q(807 downto 800) <= std_logic_vector(abs(signed(v1(807 downto 800)) - signed(v2(807 downto 800))));
  q(815 downto 808) <= std_logic_vector(abs(signed(v1(815 downto 808)) - signed(v2(815 downto 808))));
  q(823 downto 816) <= std_logic_vector(abs(signed(v1(823 downto 816)) - signed(v2(823 downto 816))));
  q(831 downto 824) <= std_logic_vector(abs(signed(v1(831 downto 824)) - signed(v2(831 downto 824))));
  q(839 downto 832) <= std_logic_vector(abs(signed(v1(839 downto 832)) - signed(v2(839 downto 832))));
  q(847 downto 840) <= std_logic_vector(abs(signed(v1(847 downto 840)) - signed(v2(847 downto 840))));
  q(855 downto 848) <= std_logic_vector(abs(signed(v1(855 downto 848)) - signed(v2(855 downto 848))));
  q(863 downto 856) <= std_logic_vector(abs(signed(v1(863 downto 856)) - signed(v2(863 downto 856))));
  q(871 downto 864) <= std_logic_vector(abs(signed(v1(871 downto 864)) - signed(v2(871 downto 864))));
  q(879 downto 872) <= std_logic_vector(abs(signed(v1(879 downto 872)) - signed(v2(879 downto 872))));
  q(887 downto 880) <= std_logic_vector(abs(signed(v1(887 downto 880)) - signed(v2(887 downto 880))));
  q(895 downto 888) <= std_logic_vector(abs(signed(v1(895 downto 888)) - signed(v2(895 downto 888))));
  q(903 downto 896) <= std_logic_vector(abs(signed(v1(903 downto 896)) - signed(v2(903 downto 896))));
  q(911 downto 904) <= std_logic_vector(abs(signed(v1(911 downto 904)) - signed(v2(911 downto 904))));
  q(919 downto 912) <= std_logic_vector(abs(signed(v1(919 downto 912)) - signed(v2(919 downto 912))));
  q(927 downto 920) <= std_logic_vector(abs(signed(v1(927 downto 920)) - signed(v2(927 downto 920))));
  q(935 downto 928) <= std_logic_vector(abs(signed(v1(935 downto 928)) - signed(v2(935 downto 928))));
  q(943 downto 936) <= std_logic_vector(abs(signed(v1(943 downto 936)) - signed(v2(943 downto 936))));
  q(951 downto 944) <= std_logic_vector(abs(signed(v1(951 downto 944)) - signed(v2(951 downto 944))));
  q(959 downto 952) <= std_logic_vector(abs(signed(v1(959 downto 952)) - signed(v2(959 downto 952))));
  q(967 downto 960) <= std_logic_vector(abs(signed(v1(967 downto 960)) - signed(v2(967 downto 960))));
  q(975 downto 968) <= std_logic_vector(abs(signed(v1(975 downto 968)) - signed(v2(975 downto 968))));
  q(983 downto 976) <= std_logic_vector(abs(signed(v1(983 downto 976)) - signed(v2(983 downto 976))));
  q(991 downto 984) <= std_logic_vector(abs(signed(v1(991 downto 984)) - signed(v2(991 downto 984))));
  q(999 downto 992) <= std_logic_vector(abs(signed(v1(999 downto 992)) - signed(v2(999 downto 992))));
  q(1007 downto 1000) <= std_logic_vector(abs(signed(v1(1007 downto 1000)) - signed(v2(1007 downto 1000))));
  q(1015 downto 1008) <= std_logic_vector(abs(signed(v1(1015 downto 1008)) - signed(v2(1015 downto 1008))));
  q(1023 downto 1016) <= std_logic_vector(abs(signed(v1(1023 downto 1016)) - signed(v2(1023 downto 1016))));
end arch;